* D:\CODE\ED - PSpice\BJT\BJT Voltage Divider\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Thu May 28 06:13:49 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
